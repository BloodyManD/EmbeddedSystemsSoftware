// niosII.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module niosII (
		input  wire [3:0]  btn_export,        //        btn.export
		input  wire        clk_100_clk,       //    clk_100.clk
		input  wire        clk_50_clk,        //     clk_50.clk
		output wire [31:0] hex_export,        //        hex.export
		output wire [7:0]  led_export,        //        led.export
		input  wire        reset_100_reset_n, //  reset_100.reset_n
		input  wire        reset_50_reset_n,  //   reset_50.reset_n
		output wire [12:0] sdram_wire_addr,   // sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,     //           .ba
		output wire        sdram_wire_cas_n,  //           .cas_n
		output wire        sdram_wire_cke,    //           .cke
		output wire        sdram_wire_cs_n,   //           .cs_n
		inout  wire [31:0] sdram_wire_dq,     //           .dq
		output wire [3:0]  sdram_wire_dqm,    //           .dqm
		output wire        sdram_wire_ras_n,  //           .ras_n
		output wire        sdram_wire_we_n    //           .we_n
	);

	wire  [31:0] cpu_data_master_readdata;                                            // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                         // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                         // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [28:0] cpu_data_master_address;                                             // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                          // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                                // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                                       // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                               // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                           // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire   [3:0] cpu_data_master_burstcount;                                          // cpu:d_burstcount -> mm_interconnect_0:cpu_data_master_burstcount
	wire  [31:0] cpu_instruction_master_readdata;                                     // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                                  // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                                      // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                         // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                                // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire   [3:0] cpu_instruction_master_burstcount;                                   // cpu:i_burstcount -> mm_interconnect_0:cpu_instruction_master_burstcount
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;              // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;           // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                 // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                      // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                       // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_performance_counter_0_control_slave_readdata;      // performance_counter_0:readdata -> mm_interconnect_0:performance_counter_0_control_slave_readdata
	wire   [3:0] mm_interconnect_0_performance_counter_0_control_slave_address;       // mm_interconnect_0:performance_counter_0_control_slave_address -> performance_counter_0:address
	wire         mm_interconnect_0_performance_counter_0_control_slave_begintransfer; // mm_interconnect_0:performance_counter_0_control_slave_begintransfer -> performance_counter_0:begintransfer
	wire         mm_interconnect_0_performance_counter_0_control_slave_write;         // mm_interconnect_0:performance_counter_0_control_slave_write -> performance_counter_0:write
	wire  [31:0] mm_interconnect_0_performance_counter_0_control_slave_writedata;     // mm_interconnect_0:performance_counter_0_control_slave_writedata -> performance_counter_0:writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;                      // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;                   // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;                   // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;                       // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                          // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;                    // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                         // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;                     // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_sdram_bridge_s0_readdata;                          // sdram_bridge:s0_readdata -> mm_interconnect_0:sdram_bridge_s0_readdata
	wire         mm_interconnect_0_sdram_bridge_s0_waitrequest;                       // sdram_bridge:s0_waitrequest -> mm_interconnect_0:sdram_bridge_s0_waitrequest
	wire         mm_interconnect_0_sdram_bridge_s0_debugaccess;                       // mm_interconnect_0:sdram_bridge_s0_debugaccess -> sdram_bridge:s0_debugaccess
	wire  [26:0] mm_interconnect_0_sdram_bridge_s0_address;                           // mm_interconnect_0:sdram_bridge_s0_address -> sdram_bridge:s0_address
	wire         mm_interconnect_0_sdram_bridge_s0_read;                              // mm_interconnect_0:sdram_bridge_s0_read -> sdram_bridge:s0_read
	wire   [3:0] mm_interconnect_0_sdram_bridge_s0_byteenable;                        // mm_interconnect_0:sdram_bridge_s0_byteenable -> sdram_bridge:s0_byteenable
	wire         mm_interconnect_0_sdram_bridge_s0_readdatavalid;                     // sdram_bridge:s0_readdatavalid -> mm_interconnect_0:sdram_bridge_s0_readdatavalid
	wire         mm_interconnect_0_sdram_bridge_s0_write;                             // mm_interconnect_0:sdram_bridge_s0_write -> sdram_bridge:s0_write
	wire  [31:0] mm_interconnect_0_sdram_bridge_s0_writedata;                         // mm_interconnect_0:sdram_bridge_s0_writedata -> sdram_bridge:s0_writedata
	wire   [4:0] mm_interconnect_0_sdram_bridge_s0_burstcount;                        // mm_interconnect_0:sdram_bridge_s0_burstcount -> sdram_bridge:s0_burstcount
	wire         mm_interconnect_0_seven_seg_s1_chipselect;                           // mm_interconnect_0:seven_seg_s1_chipselect -> seven_seg:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_s1_readdata;                             // seven_seg:readdata -> mm_interconnect_0:seven_seg_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_s1_address;                              // mm_interconnect_0:seven_seg_s1_address -> seven_seg:address
	wire         mm_interconnect_0_seven_seg_s1_write;                                // mm_interconnect_0:seven_seg_s1_write -> seven_seg:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_s1_writedata;                            // mm_interconnect_0:seven_seg_s1_writedata -> seven_seg:writedata
	wire         mm_interconnect_0_green_led_s1_chipselect;                           // mm_interconnect_0:green_led_s1_chipselect -> green_led:chipselect
	wire  [31:0] mm_interconnect_0_green_led_s1_readdata;                             // green_led:readdata -> mm_interconnect_0:green_led_s1_readdata
	wire   [1:0] mm_interconnect_0_green_led_s1_address;                              // mm_interconnect_0:green_led_s1_address -> green_led:address
	wire         mm_interconnect_0_green_led_s1_write;                                // mm_interconnect_0:green_led_s1_write -> green_led:write_n
	wire  [31:0] mm_interconnect_0_green_led_s1_writedata;                            // mm_interconnect_0:green_led_s1_writedata -> green_led:writedata
	wire         mm_interconnect_0_buttons_s1_chipselect;                             // mm_interconnect_0:buttons_s1_chipselect -> buttons:chipselect
	wire  [31:0] mm_interconnect_0_buttons_s1_readdata;                               // buttons:readdata -> mm_interconnect_0:buttons_s1_readdata
	wire   [1:0] mm_interconnect_0_buttons_s1_address;                                // mm_interconnect_0:buttons_s1_address -> buttons:address
	wire         mm_interconnect_0_buttons_s1_write;                                  // mm_interconnect_0:buttons_s1_write -> buttons:write_n
	wire  [31:0] mm_interconnect_0_buttons_s1_writedata;                              // mm_interconnect_0:buttons_s1_writedata -> buttons:writedata
	wire         mm_interconnect_0_sys_clk_timer_s1_chipselect;                       // mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_readdata;                         // sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_clk_timer_s1_address;                          // mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_0_sys_clk_timer_s1_write;                            // mm_interconnect_0:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_writedata;                        // mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire         mm_interconnect_0_instruction_tcm_s2_chipselect;                     // mm_interconnect_0:instruction_tcm_s2_chipselect -> instruction_tcm:chipselect2
	wire  [31:0] mm_interconnect_0_instruction_tcm_s2_readdata;                       // instruction_tcm:readdata2 -> mm_interconnect_0:instruction_tcm_s2_readdata
	wire  [11:0] mm_interconnect_0_instruction_tcm_s2_address;                        // mm_interconnect_0:instruction_tcm_s2_address -> instruction_tcm:address2
	wire   [3:0] mm_interconnect_0_instruction_tcm_s2_byteenable;                     // mm_interconnect_0:instruction_tcm_s2_byteenable -> instruction_tcm:byteenable2
	wire         mm_interconnect_0_instruction_tcm_s2_write;                          // mm_interconnect_0:instruction_tcm_s2_write -> instruction_tcm:write2
	wire  [31:0] mm_interconnect_0_instruction_tcm_s2_writedata;                      // mm_interconnect_0:instruction_tcm_s2_writedata -> instruction_tcm:writedata2
	wire         mm_interconnect_0_instruction_tcm_s2_clken;                          // mm_interconnect_0:instruction_tcm_s2_clken -> instruction_tcm:clken2
	wire         sdram_bridge_m0_waitrequest;                                         // mm_interconnect_1:sdram_bridge_m0_waitrequest -> sdram_bridge:m0_waitrequest
	wire  [31:0] sdram_bridge_m0_readdata;                                            // mm_interconnect_1:sdram_bridge_m0_readdata -> sdram_bridge:m0_readdata
	wire         sdram_bridge_m0_debugaccess;                                         // sdram_bridge:m0_debugaccess -> mm_interconnect_1:sdram_bridge_m0_debugaccess
	wire  [26:0] sdram_bridge_m0_address;                                             // sdram_bridge:m0_address -> mm_interconnect_1:sdram_bridge_m0_address
	wire         sdram_bridge_m0_read;                                                // sdram_bridge:m0_read -> mm_interconnect_1:sdram_bridge_m0_read
	wire   [3:0] sdram_bridge_m0_byteenable;                                          // sdram_bridge:m0_byteenable -> mm_interconnect_1:sdram_bridge_m0_byteenable
	wire         sdram_bridge_m0_readdatavalid;                                       // mm_interconnect_1:sdram_bridge_m0_readdatavalid -> sdram_bridge:m0_readdatavalid
	wire  [31:0] sdram_bridge_m0_writedata;                                           // sdram_bridge:m0_writedata -> mm_interconnect_1:sdram_bridge_m0_writedata
	wire         sdram_bridge_m0_write;                                               // sdram_bridge:m0_write -> mm_interconnect_1:sdram_bridge_m0_write
	wire   [4:0] sdram_bridge_m0_burstcount;                                          // sdram_bridge:m0_burstcount -> mm_interconnect_1:sdram_bridge_m0_burstcount
	wire         mm_interconnect_1_sdram_s1_chipselect;                               // mm_interconnect_1:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_1_sdram_s1_readdata;                                 // sdram:za_data -> mm_interconnect_1:sdram_s1_readdata
	wire         mm_interconnect_1_sdram_s1_waitrequest;                              // sdram:za_waitrequest -> mm_interconnect_1:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_1_sdram_s1_address;                                  // mm_interconnect_1:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_1_sdram_s1_read;                                     // mm_interconnect_1:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_1_sdram_s1_byteenable;                               // mm_interconnect_1:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_1_sdram_s1_readdatavalid;                            // sdram:za_valid -> mm_interconnect_1:sdram_s1_readdatavalid
	wire         mm_interconnect_1_sdram_s1_write;                                    // mm_interconnect_1:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_1_sdram_s1_writedata;                                // mm_interconnect_1:sdram_s1_writedata -> sdram:az_data
	wire  [31:0] cpu_tightly_coupled_instruction_master_0_readdata;                   // mm_interconnect_2:cpu_tightly_coupled_instruction_master_0_readdata -> cpu:itcm0_readdata
	wire  [28:0] cpu_tightly_coupled_instruction_master_0_address;                    // cpu:itcm0_address -> mm_interconnect_2:cpu_tightly_coupled_instruction_master_0_address
	wire         cpu_tightly_coupled_instruction_master_0_read;                       // cpu:itcm0_read -> mm_interconnect_2:cpu_tightly_coupled_instruction_master_0_read
	wire         cpu_tightly_coupled_instruction_master_0_clken;                      // cpu:itcm0_clken -> mm_interconnect_2:cpu_tightly_coupled_instruction_master_0_clken
	wire         mm_interconnect_2_instruction_tcm_s1_chipselect;                     // mm_interconnect_2:instruction_tcm_s1_chipselect -> instruction_tcm:chipselect
	wire  [31:0] mm_interconnect_2_instruction_tcm_s1_readdata;                       // instruction_tcm:readdata -> mm_interconnect_2:instruction_tcm_s1_readdata
	wire  [11:0] mm_interconnect_2_instruction_tcm_s1_address;                        // mm_interconnect_2:instruction_tcm_s1_address -> instruction_tcm:address
	wire   [3:0] mm_interconnect_2_instruction_tcm_s1_byteenable;                     // mm_interconnect_2:instruction_tcm_s1_byteenable -> instruction_tcm:byteenable
	wire         mm_interconnect_2_instruction_tcm_s1_write;                          // mm_interconnect_2:instruction_tcm_s1_write -> instruction_tcm:write
	wire  [31:0] mm_interconnect_2_instruction_tcm_s1_writedata;                      // mm_interconnect_2:instruction_tcm_s1_writedata -> instruction_tcm:writedata
	wire         mm_interconnect_2_instruction_tcm_s1_clken;                          // mm_interconnect_2:instruction_tcm_s1_clken -> instruction_tcm:clken
	wire         irq_mapper_receiver0_irq;                                            // sys_clk_timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                            // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                            // buttons:irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu_irq_irq;                                                         // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                                      // rst_controller:reset_out -> [buttons:reset_n, cpu:reset_n, green_led:reset_n, instruction_tcm:reset, instruction_tcm:reset2, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, mm_interconnect_2:cpu_reset_reset_bridge_in_reset_reset, performance_counter_0:reset_n, rst_translator:in_reset, sdram_bridge:s0_reset, seven_seg:reset_n, sys_clk_timer:reset_n, sysid:reset_n]
	wire         rst_controller_reset_out_reset_req;                                  // rst_controller:reset_req -> [cpu:reset_req, instruction_tcm:reset_req, instruction_tcm:reset_req2, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                                       // cpu:debug_reset_request -> [rst_controller:reset_in2, rst_controller_001:reset_in2]
	wire         rst_controller_001_reset_out_reset;                                  // rst_controller_001:reset_out -> [mm_interconnect_1:sdram_bridge_m0_reset_reset_bridge_in_reset_reset, sdram:reset_n, sdram_bridge:m0_reset]

	niosII_buttons buttons (
		.clk        (clk_50_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_buttons_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_buttons_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_buttons_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_buttons_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_buttons_s1_readdata),   //                    .readdata
		.in_port    (btn_export),                              // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                 //                 irq.irq
	);

	niosII_cpu cpu (
		.clk                                 (clk_50_clk),                                        //                                  clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                                reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                                     .reset_req
		.d_address                           (cpu_data_master_address),                           //                          data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                                     .byteenable
		.d_read                              (cpu_data_master_read),                              //                                     .read
		.d_readdata                          (cpu_data_master_readdata),                          //                                     .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                                     .waitrequest
		.d_write                             (cpu_data_master_write),                             //                                     .write
		.d_writedata                         (cpu_data_master_writedata),                         //                                     .writedata
		.d_burstcount                        (cpu_data_master_burstcount),                        //                                     .burstcount
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                                     .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                                     .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //                   instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                                     .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                                     .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                                     .waitrequest
		.i_burstcount                        (cpu_instruction_master_burstcount),                 //                                     .burstcount
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                                     .readdatavalid
		.itcm0_readdata                      (cpu_tightly_coupled_instruction_master_0_readdata), // tightly_coupled_instruction_master_0.readdata
		.itcm0_address                       (cpu_tightly_coupled_instruction_master_0_address),  //                                     .address
		.itcm0_read                          (cpu_tightly_coupled_instruction_master_0_read),     //                                     .read
		.itcm0_clken                         (cpu_tightly_coupled_instruction_master_0_clken),    //                                     .clken
		.irq                                 (cpu_irq_irq),                                       //                                  irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //                  debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //                      debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                                     .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                                     .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                                     .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                                     .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                                     .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                                     .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                                     .writedata
		.dummy_ci_port                       ()                                                   //            custom_instruction_master.readra
	);

	niosII_green_led green_led (
		.clk        (clk_50_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_green_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_green_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_green_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_green_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_green_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                                 // external_connection.export
	);

	niosII_instruction_tcm instruction_tcm (
		.clk         (clk_50_clk),                                      //   clk1.clk
		.address     (mm_interconnect_2_instruction_tcm_s1_address),    //     s1.address
		.clken       (mm_interconnect_2_instruction_tcm_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_2_instruction_tcm_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_2_instruction_tcm_s1_write),      //       .write
		.readdata    (mm_interconnect_2_instruction_tcm_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_2_instruction_tcm_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_2_instruction_tcm_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                  // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),              //       .reset_req
		.address2    (mm_interconnect_0_instruction_tcm_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_instruction_tcm_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_instruction_tcm_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_instruction_tcm_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_instruction_tcm_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_instruction_tcm_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_instruction_tcm_s2_byteenable), //       .byteenable
		.clk2        (clk_50_clk),                                      //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),                  // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),              //       .reset_req
		.freeze      (1'b0)                                             // (terminated)
	);

	niosII_jtag_uart jtag_uart (
		.clk            (clk_50_clk),                                                //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	niosII_performance_counter_0 performance_counter_0 (
		.clk           (clk_50_clk),                                                          //           clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                     //         reset.reset_n
		.address       (mm_interconnect_0_performance_counter_0_control_slave_address),       // control_slave.address
		.begintransfer (mm_interconnect_0_performance_counter_0_control_slave_begintransfer), //              .begintransfer
		.readdata      (mm_interconnect_0_performance_counter_0_control_slave_readdata),      //              .readdata
		.write         (mm_interconnect_0_performance_counter_0_control_slave_write),         //              .write
		.writedata     (mm_interconnect_0_performance_counter_0_control_slave_writedata)      //              .writedata
	);

	niosII_sdram sdram (
		.clk            (clk_100_clk),                              //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_1_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_1_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_1_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_1_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_1_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_1_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_1_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_1_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_1_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (27),
		.BURSTCOUNT_WIDTH    (5),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (32),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) sdram_bridge (
		.m0_clk           (clk_100_clk),                                     //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),              // m0_reset.reset
		.s0_clk           (clk_50_clk),                                      //   s0_clk.clk
		.s0_reset         (rst_controller_reset_out_reset),                  // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_sdram_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_sdram_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_sdram_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_sdram_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_sdram_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_sdram_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_sdram_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_sdram_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_sdram_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_sdram_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (sdram_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (sdram_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (sdram_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (sdram_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (sdram_bridge_m0_writedata),                       //         .writedata
		.m0_address       (sdram_bridge_m0_address),                         //         .address
		.m0_write         (sdram_bridge_m0_write),                           //         .write
		.m0_read          (sdram_bridge_m0_read),                            //         .read
		.m0_byteenable    (sdram_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (sdram_bridge_m0_debugaccess)                      //         .debugaccess
	);

	niosII_seven_seg seven_seg (
		.clk        (clk_50_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_s1_readdata),   //                    .readdata
		.out_port   (hex_export)                                 // external_connection.export
	);

	niosII_sys_clk_timer sys_clk_timer (
		.clk        (clk_50_clk),                                    //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                       //   irq.irq
	);

	niosII_sysid sysid (
		.clock    (clk_50_clk),                                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	niosII_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                                    (clk_50_clk),                                                          //                          clk_50_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset             (rst_controller_reset_out_reset),                                      //     cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                           (cpu_data_master_address),                                             //                     cpu_data_master.address
		.cpu_data_master_waitrequest                       (cpu_data_master_waitrequest),                                         //                                    .waitrequest
		.cpu_data_master_burstcount                        (cpu_data_master_burstcount),                                          //                                    .burstcount
		.cpu_data_master_byteenable                        (cpu_data_master_byteenable),                                          //                                    .byteenable
		.cpu_data_master_read                              (cpu_data_master_read),                                                //                                    .read
		.cpu_data_master_readdata                          (cpu_data_master_readdata),                                            //                                    .readdata
		.cpu_data_master_readdatavalid                     (cpu_data_master_readdatavalid),                                       //                                    .readdatavalid
		.cpu_data_master_write                             (cpu_data_master_write),                                               //                                    .write
		.cpu_data_master_writedata                         (cpu_data_master_writedata),                                           //                                    .writedata
		.cpu_data_master_debugaccess                       (cpu_data_master_debugaccess),                                         //                                    .debugaccess
		.cpu_instruction_master_address                    (cpu_instruction_master_address),                                      //              cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                (cpu_instruction_master_waitrequest),                                  //                                    .waitrequest
		.cpu_instruction_master_burstcount                 (cpu_instruction_master_burstcount),                                   //                                    .burstcount
		.cpu_instruction_master_read                       (cpu_instruction_master_read),                                         //                                    .read
		.cpu_instruction_master_readdata                   (cpu_instruction_master_readdata),                                     //                                    .readdata
		.cpu_instruction_master_readdatavalid              (cpu_instruction_master_readdatavalid),                                //                                    .readdatavalid
		.buttons_s1_address                                (mm_interconnect_0_buttons_s1_address),                                //                          buttons_s1.address
		.buttons_s1_write                                  (mm_interconnect_0_buttons_s1_write),                                  //                                    .write
		.buttons_s1_readdata                               (mm_interconnect_0_buttons_s1_readdata),                               //                                    .readdata
		.buttons_s1_writedata                              (mm_interconnect_0_buttons_s1_writedata),                              //                                    .writedata
		.buttons_s1_chipselect                             (mm_interconnect_0_buttons_s1_chipselect),                             //                                    .chipselect
		.cpu_debug_mem_slave_address                       (mm_interconnect_0_cpu_debug_mem_slave_address),                       //                 cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                         (mm_interconnect_0_cpu_debug_mem_slave_write),                         //                                    .write
		.cpu_debug_mem_slave_read                          (mm_interconnect_0_cpu_debug_mem_slave_read),                          //                                    .read
		.cpu_debug_mem_slave_readdata                      (mm_interconnect_0_cpu_debug_mem_slave_readdata),                      //                                    .readdata
		.cpu_debug_mem_slave_writedata                     (mm_interconnect_0_cpu_debug_mem_slave_writedata),                     //                                    .writedata
		.cpu_debug_mem_slave_byteenable                    (mm_interconnect_0_cpu_debug_mem_slave_byteenable),                    //                                    .byteenable
		.cpu_debug_mem_slave_waitrequest                   (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),                   //                                    .waitrequest
		.cpu_debug_mem_slave_debugaccess                   (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),                   //                                    .debugaccess
		.green_led_s1_address                              (mm_interconnect_0_green_led_s1_address),                              //                        green_led_s1.address
		.green_led_s1_write                                (mm_interconnect_0_green_led_s1_write),                                //                                    .write
		.green_led_s1_readdata                             (mm_interconnect_0_green_led_s1_readdata),                             //                                    .readdata
		.green_led_s1_writedata                            (mm_interconnect_0_green_led_s1_writedata),                            //                                    .writedata
		.green_led_s1_chipselect                           (mm_interconnect_0_green_led_s1_chipselect),                           //                                    .chipselect
		.instruction_tcm_s2_address                        (mm_interconnect_0_instruction_tcm_s2_address),                        //                  instruction_tcm_s2.address
		.instruction_tcm_s2_write                          (mm_interconnect_0_instruction_tcm_s2_write),                          //                                    .write
		.instruction_tcm_s2_readdata                       (mm_interconnect_0_instruction_tcm_s2_readdata),                       //                                    .readdata
		.instruction_tcm_s2_writedata                      (mm_interconnect_0_instruction_tcm_s2_writedata),                      //                                    .writedata
		.instruction_tcm_s2_byteenable                     (mm_interconnect_0_instruction_tcm_s2_byteenable),                     //                                    .byteenable
		.instruction_tcm_s2_chipselect                     (mm_interconnect_0_instruction_tcm_s2_chipselect),                     //                                    .chipselect
		.instruction_tcm_s2_clken                          (mm_interconnect_0_instruction_tcm_s2_clken),                          //                                    .clken
		.jtag_uart_avalon_jtag_slave_address               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),               //         jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                 //                                    .write
		.jtag_uart_avalon_jtag_slave_read                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                  //                                    .read
		.jtag_uart_avalon_jtag_slave_readdata              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),              //                                    .readdata
		.jtag_uart_avalon_jtag_slave_writedata             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),             //                                    .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),           //                                    .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),            //                                    .chipselect
		.performance_counter_0_control_slave_address       (mm_interconnect_0_performance_counter_0_control_slave_address),       // performance_counter_0_control_slave.address
		.performance_counter_0_control_slave_write         (mm_interconnect_0_performance_counter_0_control_slave_write),         //                                    .write
		.performance_counter_0_control_slave_readdata      (mm_interconnect_0_performance_counter_0_control_slave_readdata),      //                                    .readdata
		.performance_counter_0_control_slave_writedata     (mm_interconnect_0_performance_counter_0_control_slave_writedata),     //                                    .writedata
		.performance_counter_0_control_slave_begintransfer (mm_interconnect_0_performance_counter_0_control_slave_begintransfer), //                                    .begintransfer
		.sdram_bridge_s0_address                           (mm_interconnect_0_sdram_bridge_s0_address),                           //                     sdram_bridge_s0.address
		.sdram_bridge_s0_write                             (mm_interconnect_0_sdram_bridge_s0_write),                             //                                    .write
		.sdram_bridge_s0_read                              (mm_interconnect_0_sdram_bridge_s0_read),                              //                                    .read
		.sdram_bridge_s0_readdata                          (mm_interconnect_0_sdram_bridge_s0_readdata),                          //                                    .readdata
		.sdram_bridge_s0_writedata                         (mm_interconnect_0_sdram_bridge_s0_writedata),                         //                                    .writedata
		.sdram_bridge_s0_burstcount                        (mm_interconnect_0_sdram_bridge_s0_burstcount),                        //                                    .burstcount
		.sdram_bridge_s0_byteenable                        (mm_interconnect_0_sdram_bridge_s0_byteenable),                        //                                    .byteenable
		.sdram_bridge_s0_readdatavalid                     (mm_interconnect_0_sdram_bridge_s0_readdatavalid),                     //                                    .readdatavalid
		.sdram_bridge_s0_waitrequest                       (mm_interconnect_0_sdram_bridge_s0_waitrequest),                       //                                    .waitrequest
		.sdram_bridge_s0_debugaccess                       (mm_interconnect_0_sdram_bridge_s0_debugaccess),                       //                                    .debugaccess
		.seven_seg_s1_address                              (mm_interconnect_0_seven_seg_s1_address),                              //                        seven_seg_s1.address
		.seven_seg_s1_write                                (mm_interconnect_0_seven_seg_s1_write),                                //                                    .write
		.seven_seg_s1_readdata                             (mm_interconnect_0_seven_seg_s1_readdata),                             //                                    .readdata
		.seven_seg_s1_writedata                            (mm_interconnect_0_seven_seg_s1_writedata),                            //                                    .writedata
		.seven_seg_s1_chipselect                           (mm_interconnect_0_seven_seg_s1_chipselect),                           //                                    .chipselect
		.sys_clk_timer_s1_address                          (mm_interconnect_0_sys_clk_timer_s1_address),                          //                    sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                            (mm_interconnect_0_sys_clk_timer_s1_write),                            //                                    .write
		.sys_clk_timer_s1_readdata                         (mm_interconnect_0_sys_clk_timer_s1_readdata),                         //                                    .readdata
		.sys_clk_timer_s1_writedata                        (mm_interconnect_0_sys_clk_timer_s1_writedata),                        //                                    .writedata
		.sys_clk_timer_s1_chipselect                       (mm_interconnect_0_sys_clk_timer_s1_chipselect),                       //                                    .chipselect
		.sysid_control_slave_address                       (mm_interconnect_0_sysid_control_slave_address),                       //                 sysid_control_slave.address
		.sysid_control_slave_readdata                      (mm_interconnect_0_sysid_control_slave_readdata)                       //                                    .readdata
	);

	niosII_mm_interconnect_1 mm_interconnect_1 (
		.clk_100_clk_clk                                   (clk_100_clk),                              //                                 clk_100_clk.clk
		.sdram_bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),       // sdram_bridge_m0_reset_reset_bridge_in_reset.reset
		.sdram_bridge_m0_address                           (sdram_bridge_m0_address),                  //                             sdram_bridge_m0.address
		.sdram_bridge_m0_waitrequest                       (sdram_bridge_m0_waitrequest),              //                                            .waitrequest
		.sdram_bridge_m0_burstcount                        (sdram_bridge_m0_burstcount),               //                                            .burstcount
		.sdram_bridge_m0_byteenable                        (sdram_bridge_m0_byteenable),               //                                            .byteenable
		.sdram_bridge_m0_read                              (sdram_bridge_m0_read),                     //                                            .read
		.sdram_bridge_m0_readdata                          (sdram_bridge_m0_readdata),                 //                                            .readdata
		.sdram_bridge_m0_readdatavalid                     (sdram_bridge_m0_readdatavalid),            //                                            .readdatavalid
		.sdram_bridge_m0_write                             (sdram_bridge_m0_write),                    //                                            .write
		.sdram_bridge_m0_writedata                         (sdram_bridge_m0_writedata),                //                                            .writedata
		.sdram_bridge_m0_debugaccess                       (sdram_bridge_m0_debugaccess),              //                                            .debugaccess
		.sdram_s1_address                                  (mm_interconnect_1_sdram_s1_address),       //                                    sdram_s1.address
		.sdram_s1_write                                    (mm_interconnect_1_sdram_s1_write),         //                                            .write
		.sdram_s1_read                                     (mm_interconnect_1_sdram_s1_read),          //                                            .read
		.sdram_s1_readdata                                 (mm_interconnect_1_sdram_s1_readdata),      //                                            .readdata
		.sdram_s1_writedata                                (mm_interconnect_1_sdram_s1_writedata),     //                                            .writedata
		.sdram_s1_byteenable                               (mm_interconnect_1_sdram_s1_byteenable),    //                                            .byteenable
		.sdram_s1_readdatavalid                            (mm_interconnect_1_sdram_s1_readdatavalid), //                                            .readdatavalid
		.sdram_s1_waitrequest                              (mm_interconnect_1_sdram_s1_waitrequest),   //                                            .waitrequest
		.sdram_s1_chipselect                               (mm_interconnect_1_sdram_s1_chipselect)     //                                            .chipselect
	);

	niosII_mm_interconnect_2 mm_interconnect_2 (
		.clk_50_clk_clk                                    (clk_50_clk),                                        //                               clk_50_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset             (rst_controller_reset_out_reset),                    //          cpu_reset_reset_bridge_in_reset.reset
		.cpu_tightly_coupled_instruction_master_0_address  (cpu_tightly_coupled_instruction_master_0_address),  // cpu_tightly_coupled_instruction_master_0.address
		.cpu_tightly_coupled_instruction_master_0_read     (cpu_tightly_coupled_instruction_master_0_read),     //                                         .read
		.cpu_tightly_coupled_instruction_master_0_readdata (cpu_tightly_coupled_instruction_master_0_readdata), //                                         .readdata
		.cpu_tightly_coupled_instruction_master_0_clken    (cpu_tightly_coupled_instruction_master_0_clken),    //                                         .clken
		.instruction_tcm_s1_address                        (mm_interconnect_2_instruction_tcm_s1_address),      //                       instruction_tcm_s1.address
		.instruction_tcm_s1_write                          (mm_interconnect_2_instruction_tcm_s1_write),        //                                         .write
		.instruction_tcm_s1_readdata                       (mm_interconnect_2_instruction_tcm_s1_readdata),     //                                         .readdata
		.instruction_tcm_s1_writedata                      (mm_interconnect_2_instruction_tcm_s1_writedata),    //                                         .writedata
		.instruction_tcm_s1_byteenable                     (mm_interconnect_2_instruction_tcm_s1_byteenable),   //                                         .byteenable
		.instruction_tcm_s1_chipselect                     (mm_interconnect_2_instruction_tcm_s1_chipselect),   //                                         .chipselect
		.instruction_tcm_s1_clken                          (mm_interconnect_2_instruction_tcm_s1_clken)         //                                         .clken
	);

	niosII_irq_mapper irq_mapper (
		.clk           (clk_50_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_50_reset_n),                  // reset_in0.reset
		.reset_in1      (~reset_100_reset_n),                 // reset_in1.reset
		.reset_in2      (cpu_debug_reset_request_reset),      // reset_in2.reset
		.clk            (clk_50_clk),                         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_50_reset_n),                  // reset_in0.reset
		.reset_in1      (~reset_100_reset_n),                 // reset_in1.reset
		.reset_in2      (cpu_debug_reset_request_reset),      // reset_in2.reset
		.clk            (clk_100_clk),                        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
